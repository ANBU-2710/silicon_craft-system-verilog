interface fa_if;
  
  logic a,b,c_in;
  logic sum,c_out;
  
endinterface
